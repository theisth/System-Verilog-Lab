/*tb_lab3_g14_p2.sv
Hazirlayanlar:
Ahmet Ali Tilkicioglu
Muhammed Furkan Sarikaya
*/

`timescale 1ns/1ps
module tb_lab3_g14_p2();
logic [3:0] data;
logic [1:0] s;
logic y;
logic a;
logic b;
logic y_and;
logic y_or;
logic y_nand;
logic y_nor;
logic [7:0] data_8;
logic [2:0] s3;
logic y_8x1;
logic [15:0] data_16;
logic [3:0] s4;
logic y_16x1;

/*
mux4x1 mut0(data,s,y);
initial begin
	for (int i = 0; i < 16; i++) begin
		data = i;
		for (int j = 0; j < 4; j++) begin
			s = j;
			#10;
		end
	end 
	$stop;

end

endmodule
*/

/*
gates_mux2_1 mut0(a,b,y_and,y_or,y_nand,y_nor);
initial begin
	a = 0;	b = 0;	#10
	b = 1;		#10
	a = 1;	b = 0;	#10
	b = 1;		#10
	$stop;
end

endmodule
*/

/*
mux8x1 mut0(data_8,s3,y_8x1);
initial begin
	for (int i = 0; i < 256; i++) begin
		data_8 = i;
		for(int j = 0; j < 8; j++) begin
			s3 = j;
			#10;
		end
	end
	$stop;
end

endmodule 
*/


mux16x1 mut0(data_16,s4,y_16x1);
initial begin
	for(int i = 0; i < 65.536; i++) begin
		data_16 = i;
		for(int j = 0; j < 16; j++) begin
			s4 = j;
			#10;
		end
	end
end

endmodule


