`timescale 1ns/1ps
module tb_lab2_g14_p1_2();

logic a,b,c,d;
logic y;

lab2_g14_p1_2 mut0(a,b,c,d,y);

initial begin
	a = 0;	b = 0;	c = 0;	d = 0;	#10 //0000
	d = 1;				#10 //0001
	d = 0;	c = 1;			#10 //0010
	d = 1;				#10 //0011
	d = 0;	c = 0;	b = 1;		#10 //0100
	d = 1;				#10 //0101
	d = 0;	c = 1;			#10 //0110
	d = 1;				#10 //0111
	a = 1;	b = 0;	c = 0;	d = 0;	#10 //1000
	d = 1;				#10 //1001
	d = 0;	c = 1;			#10 //1010
	d = 1;				#10 //1011
	d = 0;	c = 0;	b = 1;		#10 //1100
	d = 1;				#10 //1101
	d = 0;	c = 1;			#10 //1110
	d = 1;				#10 //1111
	$stop;
end
endmodule