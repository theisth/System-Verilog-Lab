`timescale 1ns/1ps
module tb_deneme_1;

logic clk;
logic rst_n;
logic en;
logic [4:0] psc;
logic tick;

counter uut (
    .clk(clk),
    .rst_n(rst_n),
    .en(en),
    .psc(psc),
    .tick(tick)
);

always begin
    #5 clk = ~clk;
end

initial begin
    clk = 0;
    rst_n = 1;
    en = 0;
    psc = 5'd3;

    #10 rst_n = 0;
    #10 en = 1;

    #1000 $finish;
end

endmodule

